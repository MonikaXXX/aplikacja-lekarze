�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqK
X   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   P1q0X   P2q1X   P3q2X   P4q3X   P5q4X   P6q5etq6bX   n_features_in_q7KX
   n_outputs_q8KX   classes_q9h"h#K �q:h%�q;Rq<(KK�q=h)X   i8q>���q?Rq@(KX   <qANNNJ����J����K tqBb�C               qCtqDbX
   n_classes_qEKX   base_estimator_qFhX   estimators_qG]qH(h)�qI}qJ(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h7Kh8Kh9h"h#K �qKh%�qLRqM(KK�qNh)X   f8qO���qPRqQ(KhANNNJ����J����K tqRb�C              �?qStqTbhEcnumpy.core.multiarray
scalar
qUh@C       qV�qWRqXX   max_features_qYKX   tree_qZcsklearn.tree._tree
Tree
q[Kh"h#K �q\h%�q]Rq^(KK�q_h@�C       q`tqabK�qbRqc}qd(hKX
   node_countqeKX   nodesqfh"h#K �qgh%�qhRqi(KK�qjh)X   V56qk���qlRqm(Kh-N(X
   left_childqnX   right_childqoX   featureqpX	   thresholdqqX   impurityqrX   n_node_samplesqsX   weighted_n_node_samplesqttqu}qv(hnh)X   i8qw���qxRqy(KhANNNJ����J����K tqzbK �q{hohyK�q|hphyK�q}hqhQK�q~hrhQK �qhshyK(�q�hthQK0�q�uK8KKtq�b�Bh         
                    @�8��8��?             H@       	                    @8�Z$���?             :@                           @      �?              @                           @      �?             @������������������������       �                     �?������������������������       �                     @                           @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@������������������������       �                     6@q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KKKK�q�hQ�C�      @      F@      @      6@      @      @      �?      @      �?                      @      @      �?      @                      �?              2@              6@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       q��q�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheK	hfh"h#K �q�h%�q�Rq�(KK	�q�hm�B�                             @      �?!             H@                           @d}h���?             ,@������������������������       �                     �?                           @8�Z$���?             *@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     A@q�tq�bh�h"h#K �q�h%�q�Rq�(KK	KK�q�hQ�C�      @     �F@      @      &@      �?               @      &@       @      �?              �?       @                      $@              A@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       q��q�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheK	hfh"h#K �q�h%�q�Rq�(KK	�q�hm�B�                             @      �?             H@������������������������       �                     @                           @���7�?             F@                           @z�G�z�?             $@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     A@q�tq�bh�h"h#K �q�h%�q�Rq�(KK	KK�q�hQ�C�      @      E@      @               @      E@       @       @       @      �?              �?       @                      @              A@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       qԆq�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheKhfh"h#K �q�h%�q�Rq�(KK�q�hm�Bh                             @�q�q��?             H@                           @����X�?             ,@                           @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     @       
                     @г�wY;�?             A@       	                    @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@q�tq�bh�h"h#K �q�h%�q�Rq�(KKKK�q�hQ�C�      &@     �B@      $@      @      $@      �?              �?      $@                      @      �?     �@@      �?      @              @      �?                      <@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       q�q�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheKhfh"h#K �r   h%�r  Rr  (KK�r  hm�Bh                              @�8��8��?#             H@                           @      �?	             (@������������������������       �                      @                           @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?       
                    @������?             B@       	                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ?@r  tr  bh�h"h#K �r  h%�r  Rr  (KKKK�r	  hQ�C�      @      F@      @      "@       @              �?      "@              "@      �?              �?     �A@      �?      @      �?                      @              ?@r
  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h7Kh8Kh9h"h#K �r  h%�r  Rr  (KK�r  hQ�C              �?r  tr  bhEhUh@C       r  �r  Rr  hYKhZh[Kh"h#K �r  h%�r  Rr  (KK�r  h@�C       r  tr  bK�r  Rr  }r  (hKheKhfh"h#K �r   h%�r!  Rr"  (KK�r#  hm�Bh                             @ �q�q�?             H@                           @�q�q�?             @������������������������       �                     �?                            @      �?              @������������������������       �                     �?������������������������       �                     �?       
                    @����?�?            �F@       	                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �E@r$  tr%  bh�h"h#K �r&  h%�r'  Rr(  (KKKK�r)  hQ�C�       @      G@      �?       @              �?      �?      �?              �?      �?              �?      F@      �?      �?              �?      �?                     �E@r*  tr+  bubhhubh)�r,  }r-  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h7Kh8Kh9h"h#K �r.  h%�r/  Rr0  (KK�r1  hQ�C              �?r2  tr3  bhEhUh@C       r4  �r5  Rr6  hYKhZh[Kh"h#K �r7  h%�r8  Rr9  (KK�r:  h@�C       r;  tr<  bK�r=  Rr>  }r?  (hK heKhfh"h#K �r@  h%�rA  RrB  (KK�rC  hm�C8������������������������       �                     H@rD  trE  bh�h"h#K �rF  h%�rG  RrH  (KKKK�rI  hQ�C              H@rJ  trK  bubhhubh)�rL  }rM  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h7Kh8Kh9h"h#K �rN  h%�rO  RrP  (KK�rQ  hQ�C              �?rR  trS  bhEhUh@C       rT  �rU  RrV  hYKhZh[Kh"h#K �rW  h%�rX  RrY  (KK�rZ  h@�C       r[  tr\  bK�r]  Rr^  }r_  (hKheKhfh"h#K �r`  h%�ra  Rrb  (KK�rc  hm�B�                             @r�q��?             H@������������������������       �                     @                           @�C��2(�?             F@                           @�<ݚ�?             "@������������������������       �                     @                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?	                           @ >�֕�?            �A@
                           @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     >@rd  tre  bh�h"h#K �rf  h%�rg  Rrh  (KKKK�ri  hQ�C�       @      D@      @              @      D@       @      @              @       @      �?       @                      �?       @     �@@       @      @              @       @                      >@rj  trk  bubhhubh)�rl  }rm  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h7Kh8Kh9h"h#K �rn  h%�ro  Rrp  (KK�rq  hQ�C              �?rr  trs  bhEhUh@C       rt  �ru  Rrv  hYKhZh[Kh"h#K �rw  h%�rx  Rry  (KK�rz  h@�C       r{  tr|  bK�r}  Rr~  }r  (hKheKhfh"h#K �r�  h%�r�  Rr�  (KK�r�  hm�Bh                             @8��8���?             H@                           @      �?             @                           @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @       
                    @���N8�?             E@       	                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �C@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hQ�C�      @     �E@      @      @      @      �?      @                      �?               @       @      D@       @      �?              �?       @                     �C@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheKhfh"h#K �r�  h%�r�  Rr�  (KK�r�  hm�Bh                             @      �?             H@                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?       
                    @����?�?            �F@                           @r�q��?             @������������������������       �                      @       	                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �C@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKKK�r�  hQ�C�      @     �F@       @      �?       @                      �?      �?      F@      �?      @               @      �?      @      �?                      @             �C@r�  tr�  bubhhubehhub.